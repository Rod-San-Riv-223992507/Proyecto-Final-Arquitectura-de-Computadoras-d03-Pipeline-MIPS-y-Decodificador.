module MEM_WR(
    input clk,
    input reset,
    // Señales de control
    input reg_write_in, mem_to_reg_in,
    // Datos
    input [31:0] read_data_in,
    input [31:0] alu_result_in,
    input [4:0] write_reg_in,
    
    output reg reg_write_out, mem_to_reg_out,
    output reg [31:0] read_data_out,
    output reg [31:0] alu_result_out,
    output reg [4:0] write_reg_out
);
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            reg_write_out <= 1'b0; mem_to_reg_out <= 1'b0;
            read_data_out <= 32'b0;
            alu_result_out <= 32'b0;
            write_reg_out <= 5'b0;
        end else begin
            reg_write_out <= reg_write_in; mem_to_reg_out <= mem_to_reg_in;
            read_data_out <= read_data_in;
            alu_result_out <= alu_result_in;
            write_reg_out <= write_reg_in;
        end
    end
endmodule
